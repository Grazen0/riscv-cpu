module top_nes_bridge (
    input wire clk,
    input wire rst_n,

    output wire [7:0] led
);
endmodule
