`ifndef CPU_CSR_FILE_VH
`define CPU_CSR_FILE_VH

`define CSR_MTVEC 12'h305
`define CSR_MEPC 12'h341

`endif
