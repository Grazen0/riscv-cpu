`ifndef CPU_ALU_VH
`define CPU_ALU_VH

`define ALU_ADD 4'b0000
`define ALU_SUB 4'b1000
`define ALU_SLL 4'b0001
`define ALU_SLT 4'b0010
`define ALU_SLTU 4'b0011
`define ALU_XOR 4'b0100
`define ALU_SRL 4'b0101
`define ALU_SRA 4'b1101
`define ALU_OR 4'b0110
`define ALU_AND 4'b0111
`define ALU_PASS_A 4'b1001
`define ALU_PASS_B 4'b1010
`define ALU_AND_NOT 4'b1011

`endif
